module IM(
    input [31:0] addr,
    output [31:0] Instr
);

reg [31:0] ROM [0:4095];

wire [31:0] temp;

initial begin
    $readmemh("code.txt",ROM,0,4095);
end

assign temp = ((addr - 32'h00003000) >> 2);

assign Instr = ROM[temp];

endmodule